module core

pub struct ZOSNode {
pub mut:
	cid string // reference to circle e.g. sj4
	oid string // reference to object id in circle e.g. '3fgs'
}
