module core

pub struct ZOSClient {
pub mut:
	ref string
}
