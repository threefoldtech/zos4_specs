module cloudbox

pub struct Farmer{
pub mut:
	id string //unique id, is like key of the NFT
	
}

