module zos

pub struct ZOSClient {
pub mut:

}

pub struct Deployment {
	gid string //global id in format $cid.$oid e.g. aaa.bbb
	description string //optional, kept in circle responsible for this deployment
	
}
