module core

@[paras]
pub struct VDCSelectionArgs {
	vdcref string
}
